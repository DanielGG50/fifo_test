parameter DATA_WIDTH = 30;
parameter NUM_ELEMENTS = 16;
